parameter WORD = 32;
parameter ADDR = 16;
parameter W_IMM = 16;

