parameter WORD = 32;
parameter ADDR = 16;

