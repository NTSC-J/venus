`ifndef _params_vh_
`define _params_vh_

parameter WORD = 32;
parameter ADDR = 16;

`endif

