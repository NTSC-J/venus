/*
 * Condition Code for jump instructions
 */

`ifndef _cc_vh_
`define _cc_vh_

`define CC_ALWAYS   3'b000
`define CC_ZERO     3'b001
`define CC_POSITIVE 3'b010
`define CC_NEGATIVE 3'b011
`define CC_CARRY    3'b100
`define CC_OVERFLOW 3'b101

`endif // _cc_vh_

